module hello;
  initial $display("Hello, DeltaHDL!");
endmodule
