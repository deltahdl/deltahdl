module arithmetic;
  initial begin
    $display("%d", 2 + 3);
    $display("%d", 10 - 4);
    $display("%d", 3 * 7);
    $display("%d", 100 / 5);
  end
endmodule
